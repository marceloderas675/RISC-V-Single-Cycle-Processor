//alu to perform arithmetic and binary operations

`include "Single Cycle Processor/adder_32b"

module alu_32b 

(
    input logic [31:0] in0, 
    input logic [31:0] in1,
    output logic [31:0] out

);

endmodule