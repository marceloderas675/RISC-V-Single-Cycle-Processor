//multiplier

module Multiplier 
(
    .in0 (in0),
    .in1 (in1),
    .out (prod)
);

prod = in0 * in1;

endmodule