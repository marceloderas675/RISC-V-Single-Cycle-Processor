//register file for reading and writing

module register_file_32b 
(
    input  logic clk,
    input  logic wen,
    input  logic waddr,
    input  logic wdata,
    input  logic raddr0,
    output logic rdata0,
    input  logic raddr1,
    output logic rdata1
);

endmodule